*** SPICE deck for cell function_4_size4_2Cinv_100ps_tpdf_sim{lay} from library DDII_P1-Std_Cell_Library
*** Created on Thu Jul 02, 2020 21:06:14
*** Last revised on Wed Jul 08, 2020 23:36:52
*** Written on Wed Jul 08, 2020 23:36:57 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: function_4_size4_2Cinv_100ps_tpdf_sim{lay}
Mnmos@0 net@0 x f gnd nmos-BSIM130 L=0.14U W=1.68U AS=1.558P AD=0.195P PS=8.155U PD=2.065U
Mnmos@1 gnd y net@0 gnd nmos-BSIM130 L=0.14U W=1.68U AS=0.195P AD=0.892P PS=2.065U PD=5.53U
Mnmos@2 net@1 z gnd gnd nmos-BSIM130 L=0.14U W=1.68U AS=0.892P AD=0.195P PS=5.53U PD=2.065U
Mnmos@3 f w net@1 gnd nmos-BSIM130 L=0.14U W=1.68U AS=0.195P AD=1.558P PS=2.065U PD=8.155U
Mpmos@0 f z net@9 vdd pmos L=0.14U W=11.76U AS=3.499P AD=1.558P PS=18.235U PD=8.155U
Mpmos@3 net@9 w f vdd pmos L=0.14U W=11.76U AS=1.558P AD=3.499P PS=8.155U PD=18.235U
Mpmos@4 vdd x net@9 vdd pmos L=0.14U W=11.76U AS=3.499P AD=4.792P PS=18.235U PD=16.275U
Mpmos@5 net@9 y vdd vdd pmos L=0.14U W=11.76U AS=4.792P AD=3.499P PS=16.275U PD=18.235U

* Spice Code nodes in cell cell 'function_4_size4_2Cinv_100ps_tpdf_sim{lay}'
vdd vdd 0 dc 1.8
vx x 0 DC pulse 0 1.8 0n 100p 100p 20n 50n
cload f 0 260fF
vy y 0 dc 1.8
vw w 0 dc 0
vz z 0 dc 0
.tran 0 500n
.measure tpdf trig v(x) val=0.9 rise=1 TARG v(f) val=0.9 fall=1
.include D:\6th semester\Digital Design II\Projects\Project 1\Standard Cell Library\BSIM4_130nm.txt
.END
